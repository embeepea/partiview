89
and.cdf
ant.cdf
aps.cdf
aql.cdf
aqr.cdf
ara.cdf
ari.cdf
aur.cdf
boo.cdf
cae.cdf
cam.cdf
cap.cdf
car.cdf
cas.cdf
cen.cdf
cep.cdf
cet.cdf
cha.cdf
cir.cdf
cma.cdf
cmi.cdf
cnc.cdf
col.cdf
com.cdf
cra.cdf
crb.cdf
crt.cdf
cru.cdf
crv.cdf
cvn.cdf
cyg.cdf
del.cdf
dor.cdf
dra.cdf
equ.cdf
eri.cdf
for.cdf
gem.cdf
gru.cdf
her.cdf
hor.cdf
hya.cdf
hyi.cdf
ind.cdf
lac.cdf
leo.cdf
lep.cdf
lib.cdf
lmi.cdf
lup.cdf
lyn.cdf
lyr.cdf
men.cdf
mic.cdf
mon.cdf
mus.cdf
nor.cdf
oct.cdf
oph.cdf
ori.cdf
pav.cdf
peg.cdf
per.cdf
phe.cdf
pic.cdf
psa.cdf
psc.cdf
pup.cdf
pyx.cdf
ret.cdf
scl.cdf
sco.cdf
sct.cdf
serh.cdf
sert.cdf
sex.cdf
sge.cdf
sgr.cdf
tau.cdf
tel.cdf
tra.cdf
tri.cdf
tuc.cdf
uma.cdf
umi.cdf
vel.cdf
vir.cdf
vol.cdf
vul.cdf
